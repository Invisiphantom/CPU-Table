module Regs();
    
endmodule