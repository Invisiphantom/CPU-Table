module PCIncre(
    
);
    
endmodule